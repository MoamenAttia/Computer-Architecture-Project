library ieee;
use ieee.std_logic_1164.all;

entity testbench_decoder is
end testbench_decoder;

--architecture a_testbench_decoder of testbench_decoder is
  --  type testbench_decoder is array(0 TO 16) OF std_logic_vector(15 DOWNTO 0);
    -- signal outCases: testbench_decoder;
    -- outCases(0)  <= "0000000000000000";
    -- outCases(1)  <= "0000000000000001";
    -- outCases(2)  <= "0000000000000010";
    -- outCases(3)  <= "0000000000000100";
    -- outCases(4)  <= "0000000000001000";
    -- outCases(5)  <= "0000000000010000";
    -- outCases(6)  <= "0000000000100000";
    -- outCases(7)  <= "0000000001000000";
    -- outCases(8)  <= "0000000010000000";
    -- outCases(9)  <= "0000000100000000";
    -- outCases(10) <= "0000001000000000";
    -- outCases(11) <= "0000010000000000";
    -- outCases(12) <= "0000100000000000";
    -- outCases(13) <= "0001000000000000";
    -- outCases(14) <= "0010000000000000";
    -- outCases(15) <= "0100000000000000";
    -- outCases(16) <= "1000000000000000";
    -- begin
      -- process()
        -- begin
            
        -- end process;
  -- end a_testbench_decoder;
